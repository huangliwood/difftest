            module TOP();
                SimTop SimTop();
            endmodule
